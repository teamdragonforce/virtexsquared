`include "ARM_Constants.v"

module Decode(
	input clk,
	input [31:0] insn,
	input [31:0] inpc,
	input [31:0] incpsr,
	output reg [31:0] op0,
	output reg [31:0] op1,
	output reg [31:0] op2,
	output reg carry,

	output [3:0] read_0,
	output [3:0] read_1,
	output [3:0] read_2,
	input [31:0] rdata_0,
	input [31:0] rdata_1,
	input [31:0] rdata_2
	);

	wire [31:0] regs0, regs1, regs2, rpc;
	wire [31:0] op0_out, op1_out, op2_out;
	wire carry_out;

	/* shifter stuff */
	wire [31:0] shift_oper;
	wire [31:0] shift_res;
	wire shift_cflag_out;

	assign regs0 = (read_0 == 4'b1111) ? rpc : rdata_0;
	assign regs1 = (read_1 == 4'b1111) ? rpc : rdata_1;
	assign regs2 = rdata_2; /* use regs2 for things that cannot be r15 */

	IREALLYHATEARMSHIFT blowme(.insn(insn),
	                           .operand(regs1),
	                           .reg_amt(regs2),
	                           .cflag_in(incpsr[`CPSR_C]),
	                           .res(shift_res),
	                           .cflag_out(shift_cflag_out));

	always @(*)
		casez (insn)
		32'b????000000??????????????1001????,	/* Multiply -- must come before ALU, because it pattern matches a specific case of ALU */
//		32'b????00001???????????????1001????,	/* Multiply long */
		32'b????00010?001111????000000000000,	/* MRS (Transfer PSR to register) */
		32'b????00010?101001111100000000????,	/* MSR (Transfer register to PSR) */
		32'b????00?10?1010001111????????????,	/* MSR (Transfer register or immediate to PSR, flag bits only) */
		32'b????00010?00????????00001001????,	/* Atomic swap */
		32'b????000100101111111111110001????,	/* Branch and exchange */
		32'b????000??0??????????00001??1????,	/* Halfword transfer - register offset */
		32'b????000??1??????????00001??1????,	/* Halfword transfer - register offset */
		32'b????011????????????????????1????,	/* Undefined. I hate ARM */
		32'b????01??????????????????????????,	/* Single data transfer */
		32'b????100?????????????????????????,	/* Block data transfer */
		32'b????101?????????????????????????,	/* Branch */
		32'b????110?????????????????????????,	/* Coprocessor data transfer */
		32'b????1110???????????????????0????,	/* Coprocessor data op */
		32'b????1110???????????????????1????,	/* Coprocessor register transfer */
		32'b????1111????????????????????????:	/* SWI */
			rpc = inpc - 8;
		32'b????00??????????????????????????:	/* ALU */
			rpc = inpc - (insn[25] ? 8 : (insn[4] ? 12 : 8));
		default:				/* X everything else out */
			rpc = 32'hxxxxxxxx;
		endcase

	always @(*) begin
		read_0 = 4'hx;
		read_1 = 4'hx;
		read_2 = 4'hx;
		
		casez (insn)
		32'b????000000??????????????1001????:	/* Multiply -- must come before ALU, because it pattern matches a specific case of ALU */
		begin
			read_0 = insn[15:12]; /* Rn */
			read_1 = insn[3:0];   /* Rm */
			read_2 = insn[11:8];  /* Rs */
		end
//		32'b????00001???????????????1001????,	/* Multiply long */
//			read_0 = insn[11:8]; /* Rn */
//			read_1 = insn[3:0];   /* Rm */
//			read_2 = 4'b0;       /* anyus */
		32'b????00010?001111????000000000000:	/* MRS (Transfer PSR to register) */
		begin end
		32'b????00010?101001111100000000????,	/* MSR (Transfer register to PSR) */
		32'b????00?10?1010001111????????????:	/* MSR (Transfer register or immediate to PSR, flag bits only) */
			read_0 = insn[3:0];	/* Rm */
		32'b????00??????????????????????????:	/* ALU */
		begin
			read_0 = insn[19:16]; /* Rn */
			read_1 = insn[3:0];   /* Rm */
			read_2 = insn[11:8];  /* Rs for shift */
		end
		32'b????00010?00????????00001001????:	/* Atomic swap */
		begin
			read_0 = insn[19:16]; /* Rn */
			read_1 = insn[3:0];   /* Rm */
		end
		32'b????000100101111111111110001????:	/* Branch and exchange */
			read_0 = insn[3:0];   /* Rn */
		32'b????000??0??????????00001??1????:	/* Halfword transfer - register offset */
		begin
			read_0 = insn[19:16];
			read_1 = insn[3:0];
		end
		32'b????000??1??????????00001??1????:	/* Halfword transfer - immediate offset */
		begin
			read_0 = insn[19:16];
		end
		32'b????011????????????????????1????:	/* Undefined. I hate ARM */
		begin end
		32'b????01??????????????????????????:	/* Single data transfer */
		begin
			read_0 = insn[19:16]; /* Rn */
			read_1 = insn[3:0];   /* Rm */
		end
		32'b????100?????????????????????????:	/* Block data transfer */
			read_0 = insn[19:16];
		32'b????101?????????????????????????:	/* Branch */
		begin end
		32'b????110?????????????????????????:	/* Coprocessor data transfer */
			read_0 = insn[19:16];
		32'b????1110???????????????????0????:	/* Coprocessor data op */
		begin end
		32'b????1110???????????????????1????:	/* Coprocessor register transfer */
			read_0 = insn[15:12];
		32'b????1111????????????????????????:	/* SWI */
		begin end
		default:
			$display("Undecoded instruction");
		endcase
	end
	
	always @(*) begin
		op0_out = 32'hxxxxxxxx;
		op1_out = 32'hxxxxxxxx;
		op2_out = 32'hxxxxxxxx;
		carry_out = 1'bx;
		casez (insn)
		32'b????000000??????????????1001????: begin /* Multiply */
			op0_out = regs0;
			op1_out = regs1;
			op2_out = regs2;
		end
//		32'b????00001???????????????1001????: begin /* Multiply long */
//			op1_res = regs1;
//		end
		32'b????00010?001111????000000000000: begin /* MRS (Transfer PSR to register) */
		end
        	32'b????00010?101001111100000000????: begin /* MSR (Transfer register to PSR) */
        		op0_out = regs0;
        	end
                32'b????00?10?1010001111????????????: begin /* MSR (Transfer register or immediate to PSR, flag bits only) */
                	if(insn[25]) begin     /* the constant case */
				op0_out = ({24'b0, insn[7:0]} >> {insn[11:8], 1'b0}) | ({24'b0, insn[7:0]} << (5'b0 - {insn[11:8], 1'b0}));
			end else begin
				op0_out = regs0;
			end
                end
		32'b????00??????????????????????????: begin /* ALU */
			op0_out = regs0;
			if(insn[25]) begin     /* the constant case */
				carry_out = incpsr[`CPSR_C];
				op1_out = ({24'b0, insn[7:0]} >> {insn[11:8], 1'b0}) | ({24'b0, insn[7:0]} << (5'b0 - {insn[11:8], 1'b0}));
			end else begin
				carry_out = shift_cflag_out;
				op1_out = shift_res;
			end
		end
		32'b????00010?00????????00001001????: begin /* Atomic swap */
			op0_out = regs0;
			op1_out = regs1;
		end
		32'b????000100101111111111110001????: begin /* Branch and exchange */
			op0_out = regs0;
		end
		32'b????000??0??????????00001??1????: begin /* Halfword transfer - register offset */
			op0_out = regs0;
			op1_out = regs1;
		end
		32'b????000??1??????????00001??1????: begin /* Halfword transfer - immediate offset */
			op0_out = regs0;
			op1_out = {24'b0, insn[11:8], insn[3:0]};
		end
		32'b????011????????????????????1????: begin /* Undefined. I hate ARM */
			/* eat shit */
		end
		32'b????01??????????????????????????: begin /* Single data transfer */
			op0_out = regs0;
			if(insn[25]) begin
				op1_out = {20'b0, insn[11:0]};
				carry_out = incpsr[`CPSR_C];
			end else begin
				op1_out = shift_res;
				carry_out = shift_cflag_out;
			end
		end
		32'b????100?????????????????????????: begin /* Block data transfer */
			op0_out = regs0;
			op1_out = {16'b0, insn[15:0]};
		end
		32'b????101?????????????????????????: begin /* Branch */
			op0_out = {{6{insn[23]}}, insn[23:0], 2'b0};
		end
		32'b????110?????????????????????????: begin /* Coprocessor data transfer */
			op0_out = regs0;
			op1_out = {24'b0, insn[7:0]};
		end
		32'b????1110???????????????????0????: begin /* Coprocessor data op */
		end
		32'b????1110???????????????????1????: begin /* Coprocessor register transfer */
			op0_out = regs0;
		end
		32'b????1111????????????????????????: begin /* SWI */
		end
		default: begin end
		endcase
	end

	always @ (posedge clk) begin
		op0 <= op0_out;   /* Rn - always */
		op1 <= op1_out; /* 'operand 2' - Rm */
		op2 <= op2_out;   /* thirdedge - Rs */
		carry <= carry_out;
	end

endmodule

module IREALLYHATEARMSHIFT(
	input [31:0] insn,
	input [31:0] operand,
	input [31:0] reg_amt,
	input cflag_in,
	output [31:0] res,
	output cflag_out
);
	wire [5:0] shift_amt;
	wire rshift_cout, is_arith, is_rot;
	wire [31:0] rshift_res;

	assign shift_amt = insn[4] ? {|reg_amt[7:5], reg_amt[4:0]}     /* reg-specified shift */
	                           : {insn[11:7] == 5'b0, insn[11:7]}; /* immediate shift */

	SuckLessShifter biteme(.oper(operand),
	                       .carryin(cflag_in),
	                       .amt(shift_amt),
	                       .is_arith(is_arith),
	                       .is_rot(is_rot),
	                       .res(rshift_res),
	                       .carryout(rshift_cout));

	always @(*)
		case (insn[6:5])
		`SHIFT_LSL: begin
			/* meaningless */
			is_rot = 1'b0;
			is_arith = 1'b0;
		end
		`SHIFT_LSR: begin
			is_rot = 1'b0;
			is_arith = 1'b0;
		end
		`SHIFT_ASR: begin
			is_rot = 1'b0;
			is_arith = 1'b1;
		end
		`SHIFT_ROR: begin
			is_rot = 1'b1;
			is_arith = 1'b0;
		end
		endcase

	always @(*)
		case (insn[6:5]) /* shift type */
		`SHIFT_LSL:
			{cflag_out, res} = {cflag_in, operand} << {insn[4] & shift_amt[5], shift_amt[4:0]};
		`SHIFT_LSR: begin
			res = rshift_res;
			cflag_out = rshift_cout;
		end
		`SHIFT_ASR: begin
			res = rshift_res;
			cflag_out = rshift_cout;
		end
		`SHIFT_ROR: begin
			if(!insn[4] && shift_amt[4:0] == 5'b0) begin /* RRX x.x */
				res = {cflag_in, operand[31:1]};
				cflag_out = operand[0];
			end else begin
				res = rshift_res;
				cflag_out = rshift_cout;
			end
		end
		endcase
endmodule

module SuckLessShifter(
	input [31:0] oper,
	input carryin,
	input [5:0] amt,
	input is_arith,
	input is_rot,
	output [31:0] res,
	output carryout
);

	wire [32:0] stage1, stage2, stage3, stage4, stage5;

	wire pushbits = is_arith & oper[31];

	/* do a barrel shift */
	assign stage1 = amt[5] ? {is_rot ? oper : {32{pushbits}}, oper[31]} : {oper, carryin};
	assign stage2 = amt[4] ? {is_rot ? stage1[15:0] : {16{pushbits}}, stage1[31:16], stage1[16]} : stage1;
	assign stage3 = amt[3] ? {is_rot ? stage2[7:0] : {8{pushbits}}, stage2[31:8], stage2[8]} : stage2;
	assign stage4 = amt[2] ? {is_rot ? stage3[3:0] : {4{pushbits}}, stage3[31:4], stage3[4]} : stage3;
	assign stage5 = amt[1] ? {is_rot ? stage4[1:0] : {2{pushbits}}, stage4[31:2], stage4[2]} : stage4;
	assign {res, carryout} = amt[0] ? {is_rot ? stage4[0] : pushbits, stage5[31:1], stage5[1]} : stage5;

endmodule

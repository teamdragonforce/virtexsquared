parameter SPAM_DID_HI = 3;

parameter SPAM_ADDR_HI = 23;
parameter SPAM_ADDR_LO = 2;
parameter SPAM_DATA_HI = 31;

parameter SPAM_DID_CONSOLE = 0;
parameter SPAM_DID_LCD = 1;

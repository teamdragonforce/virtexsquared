parameter SPAM_DID_HI = 3;

parameter SPAM_ADDR_HI = 30;
parameter SPAM_ADDR_LO = 3;
parameter SPAM_DATA_HI = 31;


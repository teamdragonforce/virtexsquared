parameter DMA_SPAM_ADDR_HI = 3;
parameter NEXT_START_REG_ADDR = 4'h0;
parameter NEXT_LEN_REG_ADDR = 4'h4;
parameter COMMAND_REG_ADDR = 4'h8;
parameter FIFO_BYTES_READ_REG_ADDR = 4'hc; 

parameter COMMAND_REGISTER_HI = 1;
parameter DMA_STOP = 2'b00;
parameter DMA_TRIGGER_ONCE = 2'b01;
parameter DMA_AUTOTRIGGER = 2'b10;


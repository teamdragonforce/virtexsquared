`include "fsab_defines.vh"

/* 16 cache entries, 64-byte long cache lines */

module DCache(
	input clk,
	
	/* ARM core interface */
	input [31:0] dc__addr_3a,
	input dc__rd_req_3a,
	input dc__wr_req_3a,
	output reg dc__rw_wait_3a,
	input [31:0] dc__wr_data_3a,
	output reg [31:0] dc__rd_data_3a,

	inout valid,
	output [FSAB_REQ_HI:0] mode,
	inout [FSAB_DID_HI:0] did,
	inout [FSAB_DID_HI:0] subdid,
  	output [FSAB_ADDR_HI:0] addr,
   	output [FSAB_LEN_HI:0]  len,
   	inout [FSAB_DATA_HI:0] data,
   	output [FSAB_MASK_HI:0] mask,
        input                  credit,	


	/* bus interface */
	output wire bus_req,
	input bus_ack,
	output reg [31:0] bus_addr = 0,
	input [31:0] bus_rdata,
	output reg [31:0] bus_wdata,
	output reg bus_rd = 0,
	output reg bus_wr = 0,
	input bus_ready);
	
	/* [31 tag 10] [9 cache index 6] [5 data index 0]
	 * so the data index is 6 bits long
	 * so the cache index is 4 bits long
	 * so the tag is 22 bits long. c.c
	 */
	
	reg cache_valid [15:0];
	reg [21:0] cache_tags [15:0];
	reg [31:0] cache_data [255:0 /* {line,word} */];

	integer i;	
	initial
		for (i = 0; i < 16; i = i + 1)
		begin
			cache_valid[i[3:0]] = 0;
			cache_tags[i[3:0]] = 0;
		end
	
	wire [5:0] didx_3a = dc__addr_3a[5:0];
	wire [3:0] didx_word_3a = didx_3a[5:2];
	wire [3:0] idx_3a = dc__addr_3a[9:6];
	wire [21:0] tag_3a = dc__addr_3a[31:10];
	
	reg [31:0] prev_addr = 32'hFFFFFFFF;
	
	wire cache_hit_3a = cache_valid[idx_3a] && (cache_tags[idx_3a] == tag_3a);
	
	wire [31:0] curdata_3a = cache_data[{idx_3a,didx_word_3a}];
	always @(*) begin
		dc__rw_wait_3a = (dc__rd_req_3a && !cache_hit_3a) || (dc__wr_req_3a && (!bus_ack || !bus_ready));
		dc__rd_data_3a = curdata_3a;
		if (!dc__rw_wait_3a && dc__rd_req_3a)
			$display("DCACHE: READ COMPLETE: Addr %08x, data %08x", dc__addr_3a, dc__rd_data_3a);
	end
	
	reg [3:0] cache_fill_pos = 0;
	assign bus_req = (dc__rd_req_3a && !cache_hit_3a) || dc__wr_req_3a;
	always @(*)
	begin
		bus_rd = 0;
		bus_wr = 0;
		bus_addr = 0;
		bus_wdata = 0;
		if (dc__rd_req_3a && !cache_hit_3a && bus_ack) begin
			bus_addr = {dc__addr_3a[31:6], cache_fill_pos[3:0], 2'b00 /* reads are 32-bits */};
			bus_rd = 1;
		end else if (dc__wr_req_3a && bus_ack) begin
			$display("DCACHE: WRITE REQUEST: Addr %08x, data %08x", dc__addr_3a, dc__wr_data_3a);
			bus_addr = dc__addr_3a;
			bus_wr = 1;
			bus_wdata = dc__wr_data_3a;
		end
	end
	
	always @(posedge clk) begin
		prev_addr <= {dc__addr_3a[31:6], 6'b0};
		if (dc__rd_req_3a && (cache_fill_pos != 0) && ((prev_addr != {dc__addr_3a[31:6], 6'b0}) || cache_hit_3a))	/* If this wasn't from the same line, or we've moved on somehow, reset the fill circuitry. */
			cache_fill_pos <= 0;
		else if (dc__rd_req_3a && !cache_hit_3a && bus_ready && bus_ack) begin	/* Started the fill, and we have data. */
			$display("DCACHE: FILL: rd addr %08x; bus addr %08x; bus data %08x, bus_req %d, bus_ack %d", dc__addr_3a, bus_addr, bus_rdata, bus_req, bus_ack);
			cache_fill_pos <= cache_fill_pos + 1;
			if (cache_fill_pos == 15) begin	/* Done? */
				cache_tags[idx_3a] <= tag_3a;
				cache_valid[idx_3a] <= 1;
			end else
				cache_valid[idx_3a] <= 0;
		end
		
		/* Split this out because XST is kind of silly about this sort of thing. */
		if ((dc__rd_req_3a && !cache_hit_3a && bus_ready && bus_ack) || (dc__wr_req_3a && cache_hit_3a))
			cache_data[dc__wr_req_3a ? {idx_3a,dc__addr_3a[5:2]} : {idx_3a,cache_fill_pos}] <= dc__wr_req_3a ? dc__wr_data_3a : bus_rdata;
	end
endmodule

module Issue(
	input clk,
	input Nrst,
	
	input stall,	/* pipeline control */
	input flush,
	
	input inbubble,	/* stage inputs */
	input [31:0] insn,
	input [31:0] inpc,
	
	output reg outbubble,	/* stage outputs */
	output reg [31:0] outpc
	/* other */
	);
	
	always @(posedge clk)
	begin
		outbubble <= inbubble;
		outpc <= inpc;
	end

`ifdef COPY_PASTA_FODDER
	/* from page 2 of ARM7TDMIvE2.pdf */
	casex (insn)
	32'b????000000??????????????1001????:	/* Multiply -- must come before ALU, because it pattern matches a specific case of ALU */
//	32'b????00001???????????????1001????:	/* Multiply long */
	32'b????00010?001111????000000000000:	/* MRS (Transfer PSR to register) */
	32'b????00010?101001111100000000????:	/* MSR (Transfer register to PSR) */
	32'b????00?10?1010001111????????????:	/* MSR (Transfer register or immediate to PSR, flag bits only) */
	32'b????00??????????????????????????:	/* ALU */
	32'b????00010?00????????00001001????:	/* Atomic swap */
	32'b????000100101111111111110001????:	/* Branch */
	32'b????000??0??????????00001??1????:	/* Halfword transfer - register offset */
	32'b????000??1??????????00001??1????:	/* Halfword transfer - register offset */
	32'b????011????????????????????1????:	/* Undefined. I hate ARM */
	32'b????01??????????????????????????:	/* Single data transfer */
	32'b????100?????????????????????????:	/* Block data transfer */
	32'b????101?????????????????????????:	/* Branch */
	32'b????110?????????????????????????:	/* Coprocessor data transfer */
	32'b????1110???????????????????0????:	/* Coprocessor data op */
	32'b????1110???????????????????1????:	/* Coprocessor register transfer */
	32'b????1111????????????????????????:	/* SWI */
	default:				/* X everything else out */
	endcase
`endif

`ifdef WIP
	/* Flag setting */
	reg use_cpsr;
	reg [15:0] use_regs;
	reg def_cpsr;
	reg [15:0] def_regs;
	
	function [15:0] idxbit;
		input [3:0] r;
		idxbit = (16'b1) << r;
	endfunction
	
	wire [3:0] rn = insn[19:16];
	wire [3:0] rd = insn[15:12];
	wire [3:0] rm = insn[3:0];
	wire [3:0] cond = insn[31:28];
	
	wire [3:0] rd_mul = insn[19:16];
	wire [3:0] rn_mul = insn[15:12];
	wire [3:0] rs_mul = insn[11:8];
	
	always @(*)
		casex (insn)
		32'b????000000??????????????1001????:	/* Multiply -- must come before ALU, because it pattern matches a specific case of ALU */
		begin
			use_cpsr = `COND_MATTERS(cond);
			use_regs = (insn[21] /* accum */ ? idxbit(rn_mul) : 0) | idxbit(rs_mul) | idxbit(rm);
			def_cpsr = insn[20] /* setcc */;
			def_regs = idxbit(rd_mul);
		end
//		32'b????00001???????????????1001????:	/* Multiply long */
		32'b????00010?001111????000000000000:	/* MRS (Transfer PSR to register) */
		32'b????00010?101001111100000000????:	/* MSR (Transfer register to PSR) */
		32'b????00?10?1010001111????????????:	/* MSR (Transfer register or immediate to PSR, flag bits only) */
		32'b????00??????????????????????????:	/* ALU */
		32'b????00010?00????????00001001????:	/* Atomic swap */
		32'b????000100101111111111110001????:	/* Branch */
		32'b????000??0??????????00001??1????:	/* Halfword transfer - register offset */
		32'b????000??1??????????00001??1????:	/* Halfword transfer - register offset */
		32'b????011????????????????????1????:	/* Undefined. I hate ARM */
		32'b????01??????????????????????????:	/* Single data transfer */
		32'b????100?????????????????????????:	/* Block data transfer */
		32'b????101?????????????????????????:	/* Branch */
		32'b????110?????????????????????????:	/* Coprocessor data transfer */
		32'b????1110???????????????????0????:	/* Coprocessor data op */
		32'b????1110???????????????????1????:	/* Coprocessor register transfer */
		32'b????1111????????????????????????:	/* SWI */
		default:				/* X everything else out */
		endcase
`endif
endmodule

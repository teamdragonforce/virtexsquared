module chipscope_icon (
CONTROL0, CONTROL3, CONTROL1, CONTROL2
);
  inout [35 : 0] CONTROL0;
  inout [35 : 0] CONTROL3;
  inout [35 : 0] CONTROL1;
  inout [35 : 0] CONTROL2;
  

endmodule
